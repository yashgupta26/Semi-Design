module orgate(a,b,y);
  
  input a,b;
  output y;
  
  or g1 (y,a,b);
  
endmodule