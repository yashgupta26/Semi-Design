module tb;
  
  reg [15:0] in;
  wire [3:0] out;
  
  encoder16x4 dut (in,out);
  
  initial begin
    $monitor("in = %b;out=%b",in,out);
    in=16'b0000_0000_0000_0001; #5
    in=16'b0000_0000_0000_0010; #5
    in=16'b0000_0000_0000_0100; #5
    in=16'b0000_0000_0000_1000; #5
    in=16'b0000_0000_0001_0000; #5
    in=16'b0000_0000_0010_0000; #5
    in=16'b0000_0000_0100_0000; #5
    in=16'b0000_0000_1000_0000; #5
    in=16'b0000_0001_0000_0000; #5
    in=16'b0000_0010_0000_0000; #5
    in=16'b0000_0100_0000_0000; #5
    in=16'b0000_1000_0000_0000; #5
    in=16'b0001_0000_0000_0000; #5
    in=16'b0010_0000_0000_0000; #5
    in=16'b0100_0000_0000_0000; #5
    in=16'b1000_0000_0000_0000; #5
    $finish;
  end
  
endmodule
