module notgate(a,y);
  
  input a;
  output y;
  
  not g1 (y,a);
  
endmodule